netcdf insitu_profile_argo_1 {
dimensions:
	Location = UNLIMITED ; // (16 currently)
variables:
	int64 Location(Location) ;
		Location:suggested_chunk_dim = 10000LL ;

// global attributes:
		string :datetimeRange = "1616598060", "1616622120" ;
		string :dataProviderOrigin = "U.S. NOAA" ;
		:_ioda_layout_version = 0 ;
		string :sourceFiles = "2021032418-gdas.t18z.subpfl.tm00.bufr_d" ;
		string :source = "NCEP data tank" ;
		string :Converter = "BUFR to IODA Converter" ;
		string :_ioda_layout = "ObsGroup" ;
		string :platformLongDescription = "ARGO profiles from subpfl: temperature and salinity" ;
		string :description = "6-hrly in situ ARGO profiles" ;
		:history = "Thu Jan 30 19:31:00 2025: ncks -v MetaData/dateTime,MetaData/latitude,MetaData/longitude,MetaData/depth,MetaData/oceanBasin,MetaData/rcptdateTime,MetaData/sequenceNumber,MetaData/stationID,ObsValue/waterTemperature,ObsValue/salinity,ObsError/waterTemperature,ObsError/salinity,PreQC/waterTemperature,PreQC/salinity -d Location,3000,3015 gdas.t18z.insitu_profile_argo.2021032418.nc4 insitu_profile_argo_1.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = 0LL ;
  		string dateTime:units = "seconds since 1970-01-01T00:00:00Z" ;
  		string dateTime:long_name = "Datetime" ;
  	float depth(Location) ;
  		depth:_FillValue = 2.147484e+09f ;
  		string depth:units = "m" ;
  		string depth:long_name = "Water depth" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 3.402823e+38f ;
  		string latitude:units = "degrees_north" ;
  		latitude:valid_range = -90.f, 90.f ;
  		string latitude:long_name = "Latitude" ;
  	float longitude(Location) ;
  		longitude:_FillValue = 3.402823e+38f ;
  		string longitude:units = "degrees_east" ;
  		longitude:valid_range = -180.f, 180.f ;
  		string longitude:long_name = "Longitude" ;
  	int oceanBasin(Location) ;
  		oceanBasin:_FillValue = 999999 ;
  		string oceanBasin:long_name = "Ocean basin" ;
  	int64 rcptdateTime(Location) ;
  		rcptdateTime:_FillValue = 0LL ;
  		string rcptdateTime:units = "seconds since 1970-01-01T00:00:00Z" ;
  		string rcptdateTime:long_name = "receipt Datetime" ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = 999999 ;
  		string sequenceNumber:long_name = "Sequence Number" ;
  	int stationID(Location) ;
  		stationID:_FillValue = 2147483647 ;
  		string stationID:long_name = "Station Identification" ;
  data:

   dateTime = 1616598720, 1616598720, 1616598720, 1616598720, 1616598720, 
      1616598720, 1616598720, 1616598720, 1616598720, 1616598720, 1616598720, 
      1616598720, 1616598720, 1616598720, 1616598720, 1616598720 ;

   depth = 3, 4, 4.9, 6, 7, 8, 9, 10, 10.8, 12, 14, 16, 18.1, 20, 21.9, 24 ;

   latitude = -8.42897, -8.42897, -8.42897, -8.42897, -8.42897, -8.42897, 
      -8.42897, -8.42897, -8.42897, -8.42897, -8.42897, -8.42897, -8.42897, 
      -8.42897, -8.42897, -8.42897 ;

   longitude = -134.1183, -134.1183, -134.1183, -134.1183, -134.1183, 
      -134.1183, -134.1183, -134.1183, -134.1183, -134.1183, -134.1183, 
      -134.1183, -134.1183, -134.1183, -134.1183, -134.1183 ;

   oceanBasin = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

   rcptdateTime = 1616612820, 1616612820, 1616612820, 1616612820, 1616612820, 
      1616612820, 1616612820, 1616612820, 1616612820, 1616612820, 1616612820, 
      1616612820, 1616612820, 1616612820, 1616612820, 1616612820 ;

   sequenceNumber = 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 
      13, 13 ;

   stationID = 5905699, 5905699, 5905699, 5905699, 5905699, 5905699, 5905699, 
      5905699, 5905699, 5905699, 5905699, 5905699, 5905699, 5905699, 5905699, 
      5905699 ;
  } // group MetaData

group: ObsError {
  variables:
  	float salinity(Location) ;
  		salinity:_FillValue = 1.e+20f ;
  		string salinity:units = "psu" ;
  		string salinity:long_name = "ObsError" ;
  	float waterTemperature(Location) ;
  		waterTemperature:_FillValue = 1.e+20f ;
  		string waterTemperature:units = "degC" ;
  		string waterTemperature:long_name = "ObsError" ;
  data:

   salinity = 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
      0.01, 0.01, 0.01, 0.01, 0.01, 0.01 ;

   waterTemperature = 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 
      0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float salinity(Location) ;
  		salinity:_FillValue = 3.402823e+38f ;
  		string salinity:units = "psu" ;
  		salinity:valid_range = 0.f, 45.f ;
  		string salinity:long_name = "salinity" ;
  	float waterTemperature(Location) ;
  		waterTemperature:_FillValue = 3.402823e+38f ;
  		string waterTemperature:units = "degC" ;
  		waterTemperature:valid_range = -10.f, 50.f ;
  		string waterTemperature:long_name = "waterTemperature" ;
  data:

   salinity = 35.283, 35.284, 35.284, 35.284, 35.285, 35.283, 35.285, 35.283, 
      35.285, 35.283, 35.284, 35.285, 35.284, 35.284, 35.284, 35.284 ;

   waterTemperature = 27.70999, 27.71401, 27.71401, 27.712, 27.71099, 
      27.71099, 27.712, 27.717, 27.71301, 27.716, 27.717, 27.716, 27.71801, 
      27.71801, 27.71801, 27.71801 ;
  } // group ObsValue

group: PreQC {
  variables:
  	int salinity(Location) ;
  		salinity:_FillValue = 999999 ;
  		string salinity:long_name = "PreQC" ;
  	int waterTemperature(Location) ;
  		waterTemperature:_FillValue = 999999 ;
  		string waterTemperature:long_name = "PreQC" ;
  data:

   salinity = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

   waterTemperature = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreQC
}
